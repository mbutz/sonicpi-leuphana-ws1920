BZh91AY&SY�4� �߀Py���߰?���P^ꪪ�@�hɉ�	���0 �`�0Ú2b`b0#L1&L0H�jzD�i����C4   h�挘� ���F	� �DBd��M2a
z5<jF�4�H<���ū�YB������� $��K���h
ɡ�@���D )`�V��m���ρ[$��u:��>/���%y2�a��6a�����j��
�M'���*�(�F]���v����(w	�_()edHZ`W���|	њ�S��
ʔ��c�fZ����d��5B�6�#�e#/�(�*X%����Thn��t坒�`��؆�ȁ�r���3ͳ!��R�bw�z��1�bcca����P�ٕ�$��Yk)H��sm�7I LXAH <�)"�E��0�E��]�iby�<#:���r�?X��~?�&Lh;Z$��f� |�����#1�����y|)y|�Ww^d� �Ճ�~�C�S�D��� �u���l�9�>�9s������l=��Q�*$�Ψ��|�,��;���	JimI��Ȇ�g	���Yb���Cy%N{&v�5e0e��7�m�g�<ޗE�IF\������z���j0���0���n��_i��s$�H�B�:�>�<���Ѹm`���	%�[Dĸ�v�Ι�8r�й9ӧ��i�L���m"�^$��@@��m�>�a�H/8�� �AM��@衢��+RD9��Y�` ,���p&���딃�6�l�C5� U*BOPԢZX6�,j�7�x�:�s �"E��h��H��l�t9� �M9�; ���}�p���N���y�����#iؖ�ʏ���-l"�  wn������˿���ǐ�%0���36�4��� ��cq4���Z
�U�?�g�& s�"47��,/�k%����QҖ]o��9
I��.b���w$S�	 ��M