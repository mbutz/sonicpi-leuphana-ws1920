BZh91AY&SY�V�� I_�Py���߰?���P�y����z�h&!�4F@ �!�hɉ�	���0 �`�0�"
�(����I�6�   ��hhɉ�	���0 �`�0�$D�h��L4D��y)����26�2�kP�,x>��2�
��.Q�0Vm��6�8b���,4j�,ݨ�1����1��Pp]j�Ҟ������7A�������"����)�3���h̛9��: !K��(�6����_3�Qd*V�q�~��i7&V������>�\��b�$��Zٛ^ݖ���<�:�d0̂Úl���X�2�`��"�qaR7��<k+��ccdsoF��^��j�X����5���b��ú�L����X� aL:ǧC/a�]��=o�缋� A燨jY�m�`0�Z���\�Uc\�o��c,$Wʢ�܉��5��z^0^�}��y�w&9�Fs��̾ɖ@��K�Hx�|Y"7�����2$��I�
��^�ɱ�ۡ��0#�T%;�;	=ILS������
ǅ3�/�Bd\C��ݵq�`0J�E��]kU��:�H���}\W��Z�.��v[���Ce̞��ZR�#�Йz2&�G�+Xo�ۦ�ݿ�CD��ܵ���h�	B	.��s��$���3+�Vs�h�,Db�Q.zpe�A�p�BZS<�t:"蹌���dE*r@\P]<h����,?V� �`F��<�����E�d�����;�:��`l���	���*P�-�c�����I ��$���0mۮ�9��m����vҝ�aE( �+�,�1����g~�+"D�R�'�	c%ڙM��Z�đ��QV&#��+a�hɊ?�՚���H�kB��.�p�!�U�