BZh91AY&SY��L� J_�Py���߰?���P�┺h$Psbh0�2d��`�i���!�jA4���CML� 2144 $B@��Da���   ����a2dɑ��4�# C �"i0�Q�iSM�4�F�=&���!:	�'����d';��}�4���M�6�;3 �i�5s���RYtCG!�l���a������Uˊ��9��tim����"��ۍI�fG$�����])b��,D�@[^�?]�m��� �r�ϗ5�\>Vf^\R��[�%��\}�Q�S������e>}�3����c5��\W�O(�o:�!�R�x��*_�+R3F�=J�d�Xf6@�G24������ZYF��W�����E0`JG�%D��@e�{�^���M���^$��G?J3@?�����[�@�c��)����鐨2ʆ|H��D]`l��T �<��{���I�U��l
�6�����2�Q�%���7� ��&H�	A��(F��3$�t+dqj��2�0�=F|ʄ�P��0�iJN�Hg8��&9�Ky�[Q��tq.`���>j8
��]kQ�"y���d���̩Ka���NMA$���z�Y:�>���,��q�Mه~q���q��1���K��[~�^�#pPډ.f2Zbu�v�FH�����j� j����[I���ֈ�.c/j)C��a�p��x@l�Eޅ�!�:l���@�"����?ۙ�fEVֆH�T8���Y�&1B�04zת��a���T!�Z�c��-�����d�L���L83�O=6��}��({۱�z�c;孁"b�# �)�1����U��nX��"J(�\�W���L����:�/3�����u�%,2�2e7�]��q�)�f?��H�
���@