BZh91AY&SYdj�H �_�Py���g߰����P���wr���j�ɠ�M&�FFA����b�LFCC �#	5=MO�OI���S2C� �A�� �J��'�Mi�    �)L�O�jf���0��@ ��Lq�P
���m��]�A(?�b��![D+�bI[P���Rl*�]B�C�vԆ��d���AVTm6j�OF��ћ	�h�����9Fk�����.F�BCBFQR�m� F���κR:�(;D1㣌��6y�^���6��j|8	
��,�ЍH_�$KT�̮B�B��H�Jc�Oլ]PZGiKU�
�h��Vi������ m\cL��ll��}"�p+d�Q%(\J	��:HVhb&n����nh�p4�aV/M���{G}�z�Q+W�Z���v���6�_��fH]m��x���@�6��F��`ȷ�T��34��)��la_�=)o�`J4�nH�������n����/��BpF/�kO�E&���@��j�U~�ͱT]D�L��5�?��}���5�fD�L����qm��0�qVl7�A j�d�40S�$�9��v�HC@b�@œ��3�iyu9@����M/wXj4�Լj�M�Kj0?e�Q�{���.�u��s	Ҕ��s<�8�������i�Ęm��*P-FQ������2�$�y�S�ш��!8b�����p4���9��A�8�����3@[���At#�V�w'q�N��P2��@t�Cb=ɎVeKBv�K�ɳ�7�DkL�o�K��s��s�s�.�Xr�(�������&��YJ<T/�!8Ƹ����)*�ăB� ��5X�e�ńm4l���H�
�W) 