BZh91AY&SY
�<� H_�py��g߰?���P�=S6@�a����i�OP�4  � ��2b`b0#L1&L0H��'�z�MG�)�=OL��P ��z��2b`b0#L1&L0H�4MS�颟�Sښ��T�P22F��3Kʦ�P�����n}P���J;F
�M�6�.�ҀV��s
�Z��5�:�dCG9�^i�
Z�<�lĪk�KM������o$��\��f����2�O)�,AH@� Gq0Y;��u�[y6���I/�^/�>�\�mK�kc	8�0h����4-�{X,����ýv���1���hb9�i2�����E�XC����V�1���m�۱�k����B���0�[��!�k�`%�Q�qj�(�6�U���խl{��-����)�d\��z�8��^!�p�L��+Q�0��P1>�T)�p-�,�g(�wF.9���eH�&��5�T�p% {PFF�Lb;0`A`�F��S8�p���#�tӖ�\GQHJ\����R���_����W��;�In\��@U<�|��Q�,���w��;rC��X�'� ��]�4�kP�)������1FeH�֩�z8�<�ZB�`�9+~��(ia�S�R]M`2��&h6�'i�\c�ar%($l	#�1VU+#ubX&L��?�u1����
(�4j
B,(D%C9�r�!���R.	l�3ǫ|��g��iJ y)���څ����@��B�j%Z��]��b���4MTX��~��#�P��ǿ̍6���e��V*#	V����tQ�E�K�q�ȶ�"H$��MjH�)uM+�F���c�iUffd	��x�ʿMm70!|$Za�?��"�(Hr�R�