BZh91AY&SY634� �߀Py���g߰����P�Б��F��0�4h4���10`��`ѐ��&��D��5=L�yO#(~�� �a��a�& �4d40	�10�AѣA��dz����4�$ɴLh��
���m��YՂP~����B�D�D9�|%n��jB�0�=�hM+uHa��xwY�1A�٪�7�f�{sDт�c��/1�	�Z5��a	�$\)U���b�?Ǻ�#�.EC�og'�ɹ?���!U#��F\�&@h����5J�쀩v��L/����*W�����
�n&Ƥ������m4�=T�SN[�|��}�i�1������ ��	R�^U
c�A6�@(P�`�4@8P0����
�_3���?�k��[��P.���T`D�ï��C�	�:���4�h򼅟��XG�juMMy����>)������DL����L���y$&�}�s�l���=��E��q��s��1f<M"�	�6J}.vGɁ�ej^�욑#ɓ��^����s �\2=!������Yn)����o3�?sӂ@��$�L߬|���p����d7�Sc��Mc�Ҙ��i�a��#�h�G�ܘ��$!�N� �U>$@`�װN7�Bu�8���p�lꁥ ���	��!�eI"��NcG ��!6�Sσ���ُPH�٣���/�O��3�fA�7a��G/gFx��l��#��<Ɏ�}T�,��|�tQ�lĂ#rfَ�7bҔ20vҕ�#4|�A��W�4䞂������Ts�}�	�7�><�m4of���7������4����ńnom?�w$S�	c3J�