BZh91AY&SY�}�k NߔPyg���߰?���  P�=h�l 2i�# `F&��4� �SP�Q� P 4h4  ��DB��S#�~�I��1LF@ њ4��q�&�a22bh�A�L $�b'��44i(�ToMQ� z<�OQaE���Lo4���0�0�ԌPaF�Blmp �4�C
�Z��p�0��L�"�!A�����p����Zl߃m��~9V�+~{��8��h=s1G��e�	Zt F5�a���y~��M�ڪ����#�cf����0��G4,L%�;r/9	�v�Fa+�p('�N�e\]E(��25����"(E�8�\�FV��"��4����Y�#opυ��j��呶5�&��^��Q,- JF������(*9s�4+ml`s�/�sɦ��ǆLl�YШ�m����Ƶd�af�R�����	�u��=1=���g�;���T���Q�e���0Ps�6Q�~'��L�m�
>	s�D�ށ�2D5��Hс1&7�@������7��I�"*���|��n���!��Oi)���Aa��Q%C��^�د��8f�B��a:d���,�� g�t��e�X�w�d�Av�\I�՟s*�u"����BՊ7W#��f�u�;���Hh:�~�2Wጪ�%�7@cV��67�Z���U���:E� ���!��*�bW�$y��=�_-U�5��("QP>0������!��U��۲��
�&�A�?K7[�_j#�A�w5��sP�LL��4졩��V�aq4<�u	|�H�?�H��ڀd�Æ�����c��Èo�-�:5U��H�S¶ڰ	��FX���M0�Z�H��@"�E!��}	��d�.$6C%22r�MN㠼#[��a��{\t��օ����.�p�!D���