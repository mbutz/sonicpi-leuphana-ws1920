BZh91AY&SY���� P_�Py����߰?���P��TL�֍IM5OI�h�4hɦ� � �A�ɓ&F�L�LD"#R<�FG�����@  �`LM&L�LM2100	"&��i=�1�ii�� d�)�B���:�L΍e�B�����?�v�ؓm��8�r���Y��gc���4qD���B��՟����*Zl�����ov�R#!���d|��rV���K�r &�������*����դ�+ �k6ON��w{�;��Δ���e8t�:�Ht�vpz�P�C)A�e����6���>�RD�D�fۅ��ư��h͢Dc~��v�δ1�3��� k��լ3-\�(��5 �Re|&�{�`����Xʉch��0椸�,�;c�s�?��,��i��<} �cY�<4<�^��?���SaQvS�a�����������p%�)w�t�����ds8�`�24X�^��)���-ׇi�!�"9���Fd���m	kuS��_.��De0Ӵď�P��Dt�$ڒ�	±��_b߲�R�8��q`G^��	t^o��ؖ[5}�9Wv���9����{�X�*�-�b;B魹�CM̟2R�-)A3�PX`��-�q�MY���\�Ƙv(�-�R+U\��Iq*��1,$�u��e��cx���B�F.�pEa��e ��r�KBeέ�A��/c0j)"�7\$D$�64��H���f� �XF�vm�*���P���m�,M����s-��X�Hv�!�Ã�%�I ���PI2`�����T_a�k���؊r$��!��<ii�a\���ⴙ���.�B)E�BC��z%r-d��$Lt��d�T(30�/
)b��U�X��H�k��.�p�!����