BZh91AY&SY���� a_�Py���g߰����P~Ur�4$��蟕P��&�4�<���@� �`�2��H�&!�@h   C�0L@0	�h�h`ba�y4h51CS�ށ@����6��0(�Q�5@�|�!�qj�������āl ���;�V�0֍4��=D0T��J�H�V%�1��6(S!�M�u��17�7�K�ŵ,��R�@���CR��G͒�$u�bM0N5P�#��G�Pޖ����	�͚c�	'�w�:lR�p��� /UQbu�,��TYC,�Mj�$1N�D�����9�64~�D���ƞ&�c ��4�Kn�2l��,�<ȵ�����KRP�R��	��	1r��٬�x�e*��M3��k�r=;2�_�!�]Uy��<���O	]���g6u(��j�����& Õ-Y��d/9��;�@���Lo���[��BoG�^#`�
FP%��kHXJ'�: '<[4e���n��I�,*Ҍ��|Щ$�`�iB�py2|����t���Π�����YnA����oY�?c��5�Ip��Zy.�[���kp��TM�˸6��i�2>	�a��3�`V��pb����H�Ӛp*�d@b�װ7�Bu�������M�����K�#�qD65K��\D�4`T��*���5#f^����$��_p�KГ��A�Ga��?f����:P)[p���@v�Y4���sBŐzwϷ
4��An2�V�R�f.�R�fd�-����Na�(�2
-?*D�����rŴ�{5%Ѹ�H:o/�X���wt# �����H�
vt5�