BZh91AY&SY�� _�Py���߰?���P�rl4 M"mL�i���ha��d�@sFLL LFi�#ɀF	�jz�葓M�mMDhh@ sFLL LFi�#ɀF��ɠ&�T�hi�G��ё�=&jbр�(V�j� �$Lk���/��?�+aa�H!���eB�9�1+5v�3��|S�&#a�3��Dp�/��7�0�h��
ZM�pN0�^��������ѥ;���m��K�q����[ �K��&b"w�q_t�O�W��K�Ђ9�M~q1��x�d�P�Q�I��(t\Q�ֳ���-P�,<4���[q��#['A��~�3ǍQW,��ǐ\��I)3�CKu#E�b�U�5��k܋*�9�LcL�0ll ko�F��3\�,R�`�id-@��]tKWY�ʰ�a��JA�т�B�6!�2�dF�|��t����XW6�`s�;'LW �{B���^�����W%�6ζ�Ɓ����y	���ۍ!�^A�Fwܯҥ�)�&B�=!��$�I�Vx��$�ځS�/� <����:�R���`K���v S;�t��ר�1��� ��~����B��S(��$�h��'�*+�ɵ�O �r�(ʲ
<���h�Yk�͆���%�'xP=iڧ�|z��2�/�*�O!1vq���=p���&%��n��4�� ԇѵw-��E��a?3&�+
67� �:�����9���:�za�^s�NV��)FU3����q$%a�V�6��Xzd^��͐B[4�a(� z��#a@3Z�PF��h�]��ϻ>��:µLB�yy�Dsn ���HT���&�3�� �!�A���x"Z$B<$�����,R���,k"�  ��U΁��:�� 7�R�wD�ز����pXVM-���L�f�v:�cv'9:i`TP(%ËX�;��L!S�p���m����_ d4�����F\d�A�#�.�p�!6:$